PK   �a,W7�5i<,  *    cirkitFile.json�]mo7��+���|�7���Hb#�eq��_7�*�o$'��߯��#�L7�kT�97^ +���l�b�X���l��R__�7���zy{ys}�����e�k��Wv~�����������Og��gw�}�����O7����EnK-�,3�W"S���܋:�E^ii*ǝ�`g��x�hvNc4v	�C�U�TE�eVs#3e���,+]Q6�(+��в��ܸ�{���ʔ��r[��y�s^�K�&��)-����&�����qN���p��pI�WD~M�'���ǉ��D�	"��P�'��1��2�$�+bմ 5MD� �^Q/���D�K"�%�?!�^��$Z]Iğ$�O�'��SD�)"���?Eğ"�O��SD�)"�4��?Mğ&�O���D�i"�4��?Cğ!���g��3D�"���?Cğ!���g���D�Y"�,��?K��g���D�9��RWƱL9�3UZ��6��E����ƺF��9"t��]۰s��ZK�0���T�MM���֕0���m�]��-{������6VAh:N�FhM��}��8��0f1����U]��4���f�3��1Z��Ju�M��,��$�j�2`.�&���siD� ���yl�m�*	M�Z[0�d��2���qN�L��9n�P�1�;�rS�%��fS�L���jcD�a�jh���ŷ)�,�Ȭ�a1��˼W:+�օr��\��:���� �=������?�#+�aUa�ό���Y.k��^e����Pi-+_�\y�
.����?��/Y�5T�1%�r\CQ�1e�i���<fU��`M	�7P�\��F���
�a�i��#�P{\CQ�qE��5�󸆢�L"{��C��u�$\s�PMϒ��jyO��B��PF�	̦���Յ�0��VP�q����XA��ws(��qD��7d(���C��-�=n�P�q��vD܍$�����I<���7�x��'�o$��O��H�	��j���I<���'��I���7���'�o$�O��H
�����?#) 8~{4�m${����rQ��&�4d`0��Ņ$�[F<b��A��j�$��<�aBs��32(H���)J1F:�}Ğc�G�9N�#��4(�-7!i�W��:�]�<��"+�sYÊ��/|Bd�'���W�P�,|��u��P&�&Z�"���B�0HbQ[�4��/`Lh�����>r���L���w�@���x��7	���p��ԹF\�0��څ����$����<wd�%(?�Lb�;-�:?�F	�����H�h�wF��Fh���aq�q��E+�*`Z�'1�#�$nSN�։�L˭�������͒X1~���#x�<��D�\Ii�Ґ6Y����5�o�ت���&ɸ�$R\)>��7zy�r�F�J#F���<�y�4(iP,��4(iP,Z�N����Mcj���S�T�4(iP,ӠX�A�L�J�A�Lc�e[,ӠX�A�L�b��*�U�4(ViP�ҠX�A�J�b��*�U�4(�iP�ӠX�A�N�b��:�u�4(�iPlҠؤA�I�b��&�M�4(6iPlҠؤA�M�b��6�m�4(�iPl��ҠئA�M�bע�j�
�ڥA�K�b��n�bΘ�$�����{�-wO er�����Ql�x[����&���*��
l�x��4)�L;��ظ`+��G[�}��B��!H��il�v�nn����	�2��`��H�\Oе��,ɆUɪ�$�O�[*���V*P8G�2m�E�	�eR�u�	�L� ��9��i��<'�2��c+�H�S���y��[�<��ck���[r�@��a�H�4S�r�R&��89��I3�-UN��D�M���ts
1i <�c��mN!&��s,��)�^O�X���S�I�b��"��s,Ѕ�)ĤA�t��z:��4(�α@�T����9�:�bl�s:�]A=�Sc��W�/�R�T�[��(�#E�؊��0�zx�/�J����w0���R����w��*�}��1Ț�	ۀ,����!+/H���3���X4��1A_&�-x�/�"��`k	�����bk�Ə6��zڈ,��R�2��`K�&,&��m��!��H�^I�5o�'f���}�^I��l��2�/j�w�]M-P��?�-�+��:O"E$�"�HQI��$RL)6��D�O��D�M�^��<~y �4�i ��`��1O�b��"�N�b��"�E�4(iP,ҠX�A�L�b��2�+��2�e�4(�iP,ӠX�A�J�b��*�U"�8�U�4(ViP�ҠX�A�N�b��:�u�D�4(�iP�ӠX�A�N�b��&�M�4(6iPl�'ҠؤA�I�b��6�m�4(�iPlӠئA�MfK�b��6�]�4(viP�ҠإA��D1�@�.er��jt)���.P�KI3G��]�F�29��5��əF�ѥL�4�@�.erEA�ѥL�'��qE��ѥL;l�]ʴ���ѥL;l�]ʤ
���R&U _�6*]�F�2��5��I@�ѥL� �@�.er��jt)�s�.P�KI3G�f
]�F�2i��j	P��i�;�c�/PK &��s,�j	Ĥ��t��@-��K���|�Z1iP<�c�/PK &��s,�j	ĤA�t��@-��D�DO�X���I���|�Z1�(F�ѥLb]�F�2�O�5���`��R��e��`��R���@�.e��`���y�5���X4�@�.e:�-P�K��Ec��R&�.P�K��]\�]J��Lb]�F�2�F�5��4}�^I�jt)�+	�@�.ez%�����q?��n�������g���ٯ������U^������Ͳ��g�|���9�_���9�;s[iy�K�)�)�E��K�X�2����OnR��ghy�:�;�|��<�P2�;SZ����-�����4'o/����P2l�ղ���LѠ�2(-s��s������6m��)汌��C�)�!f�b���SBq3��Z�)2������03��=3�;#3l��~q�OO�	�M\,g��D_��GJ���*)M�h��L:;�4��[�$mKKxD������Ȼ�b���ژ#0�,;y|�6����fM�'Ȅ�Ǜ�耓��HkDj:bP��?�4����-ϲ�A&��;A��+:G{��h�ޙ�n O�fhy�9Ê�<��c#�;���M0'Џ_5�Xe�dX�X���p#��%�O��|�@?���1|����8Z��sgy��9����2��<o a�S�Fd�r�o�	vd3KygT�Qw�M�F�h�
{u���:i�{�i;�/4n�iq�y暲�@�<Kp�fO(�L�d�/�ߏ�Q�R.)��� 	{��㛎.؛��4m��,A�ٗKM\'�.�o~�����JX�:yĬՏ�y�)��K�a���Bl��9ځC���'� ��M�і�$����!1�x��H2��ح�|#������
4 ���$��� %D�g�v� ��u �8D.�l�F0g� 6l<ځC$���� �O��!�G;p�|yz�i��u�SM]���O@� y��E�j�Ve�EK�A���(h�/	�s�ٜ��T������!8D��lCp�PK�8$V@̦�B��F ƞo��,� �)$�rp0St� l�)V�#b��T9n�lJR�B[R�W�=�V���� �,s�RR����0Ժ����g�!�V��ۣC$��{@�����Z�C\�������="/�S��uX	z@,�J�bU1���J�pz� ���lK��N�(C��;!Yul��]�PV��D��{�}U!f�Q�9[�4?��"�.$����<�G���O��`�X�:�F	[�:[�e���԰խ�� �\�N��u=%=1�b�#8H�Ô->@��li��޾������!*��x��䂃���ԌG�WJ��� :�\�p�5�v���)Nd�qU��N�=X�`�.��x��q;p�(՜#p�0�$|���41ځ�\8A=��� b58�m�1���bK�G�d�8�n}jr	�Ikx�,�/~F#�Qŧm�&̘t���e�]zY�1�l/���q���I�s�9O8r�J��9����\ì���M��5%�
��b�= ޯ�d�8�5U�f�z��qw���SK����M� ��͗�t�艆���e�������.��Ϟ��~�4�.�n.>_Vg��l��!_ ˉ���>}̶���2S=q�V��'�L����S�FF+���W.�U��
�Sqȩ@�T$
*�pR�(�H}c�)�9ѷ��R�$�8T�
*N���SIũ$��T�J�ŔT�)�H�T$J*%���DEE��"QQ���HTT$**���DEE��"QS���H�T$j*5���DME��"QS�h�H4T$*���DCE��"�P�h�H4T$Z*-���DKE��"�R�h�*-���D��1�H�0N��
LG��h���Fp�:,1�h�(@�}a�(q#fy16h�<��FȑI=q�,�����"/]��=2i�7�����(�ם2�`к3�� �~��-؛⪉����-C�6���#��u�č�A\�|��?�v8����������J����(�x#�;�^�
_�Q1�B^쪏�*gd�pW��G&w�����G\d���A�X���A�X~� �"p�'�����z�}WDT��c/#
�"q�'�l�H;��	�"QP�8v�@E��a<�FP�FE��a<N yY�"q�0'��ı�x�7D��jcg�د�`]QdQKO�ä؈�n�^�"�?��E�-=���;��N� *�x� a������ಳ�@G��E�1S���F������k(�t��ǂ��j4t�#n,x��A�FkJP�FЁ�R����`#�G�!�bI�f�n���-佛��!/2E[ULQ��"��[d0�c��({$�7��`��\�1֛C�[��?���.�P�oC%�����g���&x\a����� �o(fk����n{*���턴ǘ<��@�~�8D+;p���G�5�"p��!�2p��!��8d���C8ڏ����
�}����
*p���G{wF[����}����:p��a�	&p���~�Ǵ�8L�0��-�moIi�5`�6p����dc�m��.p����E�N�}<?Ü0�O&���퉈�5ġ��R1���T�ٱ}���07��{x͏A��fl��?�f@���#��p�P�t�
Yj�\���a��+T���s��%�e��I�c������[A��� ��̭�D�x��0W�8�@��F"yS�&��*����@Y����k���,���&�.i��ko��v�d��yeW��Rqi3YV0X�dhUg^���g��d�����5��V0���Ƹ�Jź3y�d�l{���~0肑���7uλ7*�a�����\V5��:c0�+�TkC�~�Jp�d`,a��`�u��³B��Ȼ�A�v�,�,t������2w@]7%��I������x�+&�)Z����y�IS�L�p@k�2�yÝT`��Ժ��Օ � xк40�M^
P~o:��)뺔0�����s�0��R�Hƚ�
X`�J�7F��"oL��`k�v^w��^y[����e(K�(�5���H[���(�*]�$1Ze\VxP-axYX�E#�9�kU�(� �6��LV�KU1&|�OX��� #'`��7�"dZ�5(4�*$緭U��Pw��ʺQ0���u�+�Z��K}^�P��]�.:����?���}0r���TCʥ�*zd������t�3g(3G��=~�H��g�p{eJ|�?�62���LO�3.ҙ�|�����!>X�댌t�/�u�S@C��R3ʹEt�_Lɩ�d��E����v��t�W��:sHqk[�31���^gb�� ��z���T�כ�>�z�W������U^�W���Q�����{Z�yd�G���v�l�����#�=�G�{$��x������?b�#�{��m�~c|=�?|��7��;��%_�6�7_w~�	˯�.�e�W�M��..������ۻ�#�+Y2�2f�^� ���3�L:�sf+�.��k�?yqU7w��7۷_�wa��{���˛O���n��?��p���[^^���:�9������_}��o�Fj?__B#g���O7���~	rϞ7��mo������U}��e���/�uu��^ F����3l��>/��X6�6z��A,AO�+�nn/�.o`~��,�~�Bq�qi�?���6��5�8�|"%����{-xV�c��uŹw���vy}{�_�+��������._�쬺�5LEy�,��n>�g��3a��o�S�T~��N���~A�s,<0����E��_�����m<Gq��A&���m���	�v�O�<#2Gf��8w#|f�O����V�^l�)��}O������(����(������&�1�+�>QQ�Q�Y����cO��=1Qk��ܫa2�1#��A�	�m���d�u���F23 `��w�Imk��x$ն�l<�q.�b��~o=�j�U�gz�O��m<>��os��w�>��ŹL�K�����g2�&v����x�A;խ=C3�=�����Lw��fz�hx��g�3�=�����Lw��f�{48ӫg�3�z48ӫG�3�z��\�������z84�������uy���suy�C��]�H|�O���|�-�p�	8��>�����urO���s�m7��l���4��Ӧ�[�������2Ls#3�|8,��������tQ��(O��C��`O�����Y�Z+��/�+M�z������L�6��ذ�jy�W�:�a��70��¸��®� ��'*+y�!����~2�ɚ�ՎW�m>�ZP��h��i +�[*5k�<Q�V��=�M�� X{f�<,?�h����b7����!�Yj�g��MF��l�e�*ƛ��@���� �6�ﳣ�o��Ld_��O�&��yy�~�%��Xgy�=װ�4�	�mJ��,3�Bb�
�1y�⦨�F�ڋ0�P�h�b� h�e����0)��p�� x&NK�^,�ni���� �T'�SA�Fzc:S	Mj��Y�k�9��U��!��>�} Z������������5�;��yT�
��ǵ�϶���M�`�¥�CH�]<EF���-�"bBk-⻿�`o� �mg�I������]�g��7`�g�p�)p�ͫgo߼����z��ts�//�~ې}��{��ć��(b�:?k�.?�\���^�������}�-�����sy���zysu��M�٥yx�4��~`�)/��|��5�}3|T|8�����F�WJ9���������A����&�E%mn2o>�
/�}W�:ֽmӣ�Y8넲R��3��rB3��Gi'�*��>$�*S����!�#lUX�kP���n�i���і��m)���b���B�j�l�9�������ώ.���c�E�7�ϗw�^_W��Ij,dJ��Px&�vxLo���2e�3]K�T[)2]��l�����Y��u��dP�G&��=o>���:�H�� ��S��ĕ�+Ѳݩy�6lc�I���5@��7j:`��3�/[�gQk��L�� 6Q9+3�����J�P�����'T�η~Z{»�v�����fx��;>]�BÃ�G���0��8���}��n�ywܬ7��<��5W|M�:*�3_�.�9���d]��, �g{0p�aڵ���DG�2|e��y��&DT�.��x�Lp�p�qݞ�l��5^΃#Z S��&UK�����aTt�tҒ�q.��4�h���=�&��G��f�4����@k3Z��F��A��Z���D�A�I�[���� ��+�u}r i��VH�6�n B�\j�BZ�=H���֡E������-���	�P���L���yWm�����0������#����P��̦΁�.�tEVrjq,�;X�97 ��s�*
E�|�k�H��a��~Ѧ[��ʍgBv���3���c��:$�wN����LD\���!����2����_e����7o�z� �}~�����ߞ��L�]���+�;#�̹�����Ă�%��!ԡeB�.��P�ה�f��U#{!`L2��Rs�Cb�r۾3�v�7��d��x��<"��c<��xd�C[��[���#i�Lz��:H��U�(�����x���6��$�w��`�8W��֏��#�V׫��>п�lPs,�P+}��n��_�O68T}�����V�jh��TCh�S­O6��>� ��dCӣԸ>Ր����4�O5d1�TC�O5h�zd������7Ιb�����eZ1#�}pf6ܲ�i^�*��V�gy�������8Ꞿtѫl�v���-��+m��q�hsg �Ȭ��E��@��k��' ��������/����B-l��d��د���V^3 ��bw���yi2fj��Z���������]�,/��� b��0�FѺ�BƠ�*drt����q�p��k�';2�7�&�v8�1��+N0�|���v��a7.l�B���	�*v��[��	�Q����P�`�֞l���.�87�S��I0�l�yx������go�y�����tP|ȃb�U��΃�Τv6x� ~VJ/���9*F݅4�Q�c���ó/O�x�Ń�b(�4�ڐ˝e4|�8�F��ʩ���l�	�b�ᚋ�}������񤏇]�^X'<oVL8��fa����9oOdi
����i)�>��I����5�͡���l8��F.3Fh���Պ���{3��6~���g�����IO�xH]̌�iBv�U<V��B G��b�2:�s7�S���^}����/�{������?)�I)��:\A���ʅ�h8R�f!C��Q�1饥*%��'��߿z���'�<��U��E�5���i�|8v��
2�9w�+�N�.\B:���o^��3wRƓ2R�S��F�q$�9�-h���Z��>+�OI��ճw��{��4�����j�S�J:X��]�(�tR�.RҽU�gC��:�+#?��I�2�, ���R�2h����� �UJF.G}��ɩ�8��I��r���Q2��T<�JᝲΓ�D�g���"ʓ"��hϕ��pυ3�	m���]�'��������Z�uś*�\�s��-��mF�2�-G�)!꓍OH	�v���VMȼ�S�9��9h�BX&`�R��~��������U'5<�����څ ͑6�F������{����{r6*�K�OI	O�Z	]�&�=�`e
�Z�N�9��"�W�������g�������Oǈ'�<p�wr��1NK�g��?PJ�`M4Z[/U#�Zպ�&�E��f�.:��й�	����}����)�I����1Z*�t��s��N��eN0A/`��j[�̉ڇ`p;�3���<�J�'���Cē&X�_�A��w��ܹP?�C��ËF���RdUa@K�u��4��s_9�bQ��E A��w7 ���
/��o�5��ۯ���Oa�\����a-��n/�	RqV���������� l��?��W��O~����~����0��̿ {��p��C@��
����X�|	�v��j=�S�+a�u5*
��ӊZ濾K�5��*]�>�\����~je���Ç���7����]kuo�_����q�g�9���>��k�8_�Y���Y.+ރl�.���k�T۟๧��V� ��?>���$�s�;
����qa�^z�0��.��9��Qt�!�":�0�,?�5ۣkG�Y�����)�%���AH���a�#h��{9܁�ƬMH��As��G��>};*8�/��ؾN66�8�#"q1�?0�];��лN��2��X��Џ�C!Yb�嵭Sn�T:����5�j2�v��+��0,�0��؄7���#�#0�%�jO�Т��=�v\��n�֗��)�WYX�7g�k��bێ��
�O���ql�];*h������D��cȎ �폂�}�vT�x�:b��GuDd`�hq`�vd�k�ÿ������<w,��`I�jE�cH�a�w�t�0�.�j{t�=z�'��.�S�#S|P�d�
I�e�>�l���d���TÀ�Z���t���c����c������әG�v��&�؟(����0����zb>֋����R�̚�	�l��"Z�B9_k.L�4���?��퉟���b���Q��$bB�/�?�G,Bֆ�E$����h|�������Ţ���l�KV����6h���Zg�v�i���&�܉-a�����-l��� �7T����1���[�`�)��*m��ځ���Ym��s!,S�>1�=�� ��{ ��)�퐙�~Y�Zud�C�UXw������C�,"Qv�8�ܣkGF�vT4j"wȆ�d�PC��y��D%���X��Cx��q���<E1�!�yt��ƒ!�x�&%�$Ϊa|�=�!{tc��b�Ƕ�v��Lۈ�&C&��߽kO���+���∘I��i��!�gǛ�{��O���o�q��h*� {��g������@��'�Z�gG�b���n�KƇbM;��>U���H����2���C�,��3�VJ�<�F����������5������;���]5��P�1d�;�k�$�T����T�N�ڨX�6|�Y�EQn��=����|dtѵǴζ���o�J�kѶ����;�'}�8���]K��ެ�,�=�a0�bzt�5G��;���gǃ�Z*k����,�]��,U����4�"�TrkߓJm+�Ƈ����oiR�#�FL�K�+�߈�ݾ�w;ɢ�Ļ2������bǺ�VI�\5�"������w��6�K�Md��#��y=��T;]I3v.e5E�Sv:gw��틠m�0��m��@,�ۑU4����]d�O�X$�PE'���K��ڣo ��=jE��nǩ�e17h7�h��˫�7ͷ�]��̯nϞ�ܶ�\����ͯ?�W_�������6���?���?PK
   �a,W7�5i<,  *                  cirkitFile.jsonPK      =   i,    